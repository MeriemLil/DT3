//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// sva_bindings.svh: SVA assertion module bindings for RTL simulation and formal verification.
//
// - The macro 'RTL_SIM' is defined in the RTL simulation script.
// - The macro 'design_top_is_*' is defined in the RTL simulation script based on
//   the value of the DESIGN_NAME TCL variable.
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

// This macro is defined in project-file include file audioport.svh

`ifdef INCLUDE_ASSERTIONS

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// SECTION 1: Bindings for RTL simulation.
//
//            - Hierarchical paths of instances begin from testbench module.
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef RTL_SIM

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  1.1. control_unit
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_control_unit

//       Example: Binding an assertion module to all instances of a design module
//
//       .------------------------------------------- Name of module bound to (design module)
//       |           .------------------------------- Name of module to be bound (assertion module)
//       |           |                   .----------- Instance name of module to be bound (assertion module)
//       |           |                   |
//       V           V                   V
bind control_unit control_unit_svamod CHECKER_MODULE (.*);
`endif


/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  1.2. dsp_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_dsp_unit
bind dsp_unit dsp_unit_svamod CHECKER_MODULE (.*);
`endif

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  1.3. cdc_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_cdc_unit
bind cdc_unit cdc_unit_svamod CHECKER_MODULE (.*);
`endif
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  1.4. i2s_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_i2s_unit
bind i2s_unit i2s_unit_svamod CHECKER_MODULE (.state_r_port(state_r), .*);
`endif

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  1.5. audioport
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_audioport
bind audioport audioport_svamod CHECKER_MODULE (.*);
bind control_unit control_unit_svamod CHECKER_MODULE (.*);
bind dsp_unit dsp_unit_svamod CHECKER_MODULE (.*);
bind cdc_unit cdc_unit_svamod CHECKER_MODULE (.*);
`ifndef CDS_TOOL_DEFINE
bind i2s_unit i2s_unit_svamod CHECKER_MODULE (.state_r_port(state_r), .*);
`endif
`endif


`endif //  `ifdef RTL_SIM


//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// SECTION 2: Bindings for formal verification.
//
//            - Hierarchical paths of instances begin from top module.
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifdef RTL_VERIF

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  2.1. control_unit
//
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_control_unit
bind control_unit control_unit_svamod CHECKER_MODULE (.*);
`endif


`ifdef design_top_is_bus_interface
bind bus_interface bus_interface_svamod CHECKER_MODULE (.*);
`endif

`ifdef design_top_is_cregs
bind cregs cregs_svamod CHECKER_MODULE (.*);
`endif

`ifdef design_top_is_abuf
bind abuf abuf_svamod CHECKER_MODULE (.*);
`endif


/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  2.2. dsp_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_dsp_unit
bind dsp_unit dsp_unit_svamod CHECKER_MODULE (.*);
`endif

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  2.3. cdc_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_cdc_unit
bind cdc_unit cdc_unit_svamod CHECKER_MODULE (.*);
`endif
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  2.4. i2s_unit
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_i2s_unit
bind i2s_unit i2s_unit_svamod CHECKER_MODULE (.state_r_port(state_r), .*);
`endif

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//  2.5. audioport
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef design_top_is_audioport
bind audioport audioport_svamod CHECKER_MODULE (.*);
bind control_unit control_unit_svamod CHECKER_MODULE (.*);
bind dsp_unit dsp_unit_svamod CHECKER_MODULE (.*);
bind cdc_unit cdc_unit_svamod CHECKER_MODULE (.*);
`ifndef CDS_TOOL_DEFINE
bind i2s_unit i2s_unit_svamod CHECKER_MODULE (.state_r_port(state_r), .*);
`endif
`endif

`endif


`endif
