`include "audioport.svh"

import audioport_pkg::*;
